--------------------------------------------------------------------------------
-- Create Date:    15:24:38 11/10/05
-- Design Name:    
-- Module Name:    search - Behavioral
-- Project Name:   Deflate
-- Target Device:  
-- Dependencies: Hashchain.vhdl
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- Slightly modified approach to use a hash search
-- Instead of searching a chain of hashes a table of the hashes generated by the
-- minimum length chains is maintained
--------------------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

--Function to find the log of a number 
--Is used to convert the addresses
package mat is
	 function log2(v: in natural) return natural;
end package mat;

--Function definition
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;


package body mat is

function log2(v: in natural) return natural is
	variable n: natural;
	variable logn: natural;
begin
	n := 1;
	for i in 0 to 128 loop
		logn := i;
		exit when (n>=v);
		n := n * 2;
	end loop;
	return logn;
end function log2;
end package body mat;
--End of the package



library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use work.mat.all;

entity stream_search is
	Generic 
	      (Length_of_Table : natural :=	32768;            -- Number of locations in the hash table default = 32k table
			 Hash_Width      : natural := 32;	 				-- Number of bits in the hash
			 Data_Width      : natural := 8 					-- Data bus width			 )
			 );
	Port
	      (
			Table_Start      : in    std_logic_vector ( log2(Length_of_Table) downto 0);   -- Starting Address of the data table
			Table_End        : in    std_logic_vector ( log2(Length_of_Table) downto 0);	 -- Ending address of the table
			Hash_key         : in    std_logic_vector ( (Hash_Width -1) downto 0);			 -- Accept a 32 bit hash input	
			Hash_inout		  : inout std_logic_vector ( (Data_Width -1) downto 0);			 -- Hash key read/write to be stored
			Data_in			  : in    std_logic_vector ( (Data_Width -1) downto 0);     	 -- Data input from byte stream
			Clock,						 																       -- Clock input	
			Output_E			  : in    bit;																	 -- Enable/~Tristate output
			Table_Match      : in    std_logic_vector ( log2(Length_of_Table) downto 0);   -- Address at which the match was found
			Match				  , 						  														 -- when 1 hash key generated matches hash from table 
			Write_Hash		  : out   bit																	 -- no match read the next byte from memory
			);
end stream_search;
--The search is a one to one search of the table
--The hash keys are stored FIFO unsorted in the table.
--it is the easiest method and needs to be changed to a sorted store-search.
architecture one_to_one of stream_search is
component Hash1
          Port ( 
			  Hash_o   : out std_logic_vector (Hash_Width - 1 downto 0);     -- Hash value of previous data
           Data_in  : in  std_logic_vector (Data_Width-1 downto 0);       -- Data input from byte stream
			  Clock,													                    -- Clock
			  Reset,													                    -- Reset
			  Output_E : in  bit		                     						  -- Output Enable
           );
end component;

begin


end one_to_one;
